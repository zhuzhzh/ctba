//
// Created by         : Harris Zhu
// Filename           : hw_top.sv
// Author             : Harris Zhu
// Created On         : 2016-11-15 20:35
// Last Modified      : 
// Update Count       : 2016-11-15 20:35
// Tags               :  
// Description        : 
// Conclusion         : 
//                      
//=======================================================================

module hw_top;

memBFM u_membfm();
dut u_dut();

clkgen u_clkgen();

endmodule
